`define LEVELS $clog2(FFT_SIZE)
`define BYTE_COUNT $clog2(DATA_WIDTH)
`define ADDR_WIDTH $clog2(FFT_SIZE)
`define NUM_TWIDDLES FFT_SIZE/2
