package axis_master_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "axis_trans.sv"
    `include "axis_master_driver.sv"
    `include "axis_master_seq.sv"
    `include "axis_master_agent.sv"

endpackage
