`define LEVELS $clog2(FFT_SIZE)
`define BYTE_COUNT DATA_WIDTH/8
`define ADDR_WIDTH $clog2(FFT_SIZE)
`define NUM_TWIDDLES FFT_SIZE/2
