`define LEVELS $clog2(FFT_SIZE)
`define DATA_WIDTH 2*(SAMPLE_WIDTH + $clog2(FFT_SIZE)/2)
`define IN_AXI_WIDTH SAMPLE_WIDTH
`define IN_BYTE_COUNT `IN_AXI_WIDTH/8
`define OUT_AXI_WIDTH (1 << $clog2(`DATA_WIDTH))
`define OUT_BYTE_COUNT `OUT_AXI_WIDTH/8
`define ADDR_WIDTH $clog2(FFT_SIZE)
`define NUM_TWIDDLES FFT_SIZE/2
`define TWIDDLE_WIDTH 50
