package fft_pkg;

    import uvm_pkg::*;
    import axis_master_pkg::*;
    import axis_slave_pkg::*;
    import fft_ctrl_pkg::*;

    `include "../../sources_1/new/fft_defs.vh"
    `include "uvm_macros.svh"

    `include "mem_mux/mem_mux_seq_item.sv"
    `include "mem_mux/mem_mux_monitor.sv"
    `include "mem_mux/mem_mux_scoreboard.sv"
    `include "fft_env.sv"
    `include "fft_test.sv"

endpackage
