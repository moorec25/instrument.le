package axis_slave_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "axis_slave_trans.sv"
    `include "axis_slave_monitor.sv"
    `include "axis_slave_scoreboard.sv"

endpackage
