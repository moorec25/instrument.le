class fft_ctrl_trans_t extends uvm_sequence_item;

    logic fft_start;
    
    `uvm_object_utils(fft_ctrl_trans_t);

    function new(string name = "fft_ctrl_trans_t");
        super.new(name);
    endfunction

    
endclass

