interface fft_ctrl_if_t;
    logic clk;
    logic reset;
    logic fft_go;
    logic fft_busy;
endinterface
