package fft_ctrl_pkg;
   
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "fft_ctrl_driver.sv"
    `include "fft_ctrl_seq.sv"
    `include "fft_ctrl_agent.sv"

endpackage
